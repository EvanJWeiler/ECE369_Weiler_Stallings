`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  1
// Module - InstructionMemory.v
// Description - 32-Bit wide instruction memory.
//
// INPUT:-
// Address: 32-Bit address input port.
//
// OUTPUT:-
// Instruction: 32-Bit output port.
//
// FUNCTIONALITY:-
// Similar to the DataMemory, this module should also be byte-addressed
// (i.e., ignore bits 0 and 1 of 'Address'). All of the instructions will be 
// hard-coded into the instruction memory, so there is no need to write to the 
// InstructionMemory.  The contents of the InstructionMemory is the machine 
// language program to be run on your MIPS processor.
//
//
//we will store the machine code for a code written in C later. for now initialize 
//each entry to be its index * 4 (memory[i] = i * 4;)
//all you need to do is give an address as input and read the contents of the 
//address on your output port. 
// 
//Using a 32bit address you will index into the memory, output the contents of that specific 
//address. for data memory we are using 1K word of storage space. for the instruction memory 
//you may assume smaller size for practical purpose. you can use 128 words as the size and 
//hardcode the values.  in this case you need 7 bits to index into the memory. 
//
//be careful with the least two significant bits of the 32bit address. those help us index 
//into one of the 4 bytes in a word. therefore you will need to use bit [8-2] of the input address. 


////////////////////////////////////////////////////////////////////////////////

module InstructionMemory(Address, Instruction); 

    input [31:0]Address;        // Input Address 

    output reg [31:0]Instruction;    // Instruction at memory location Address
	
	reg [31:0]memory [0:511];  
    
    /* Please fill in the implementation here */
	initial begin
	//$readmemh ("vbsme_small_stripped.mem", memory);
	//$readmemh ("vbsme_1_stripped.mem", memory);
	//$readmemh ("test5_stripped.mem", memory);
	//$readmemh ("test4_stripped.mem", memory);
	$readmemh ("Instruction_memory.mem", memory);
	//begin forwarding testing
	 /* memory[0] = 32'b00100000000100000000000000000001; //	main:	addi	$s0, $zero, 1 (s0 = 1)
      memory[1] = 32'b00100000000100010000000000000001; //        addi    $s1, $zero, 1 (s1 = 1)
      memory[2] = 32'b00000010000100011000000000100100; //        and    $s0, $s0, $s1 (s0 = 1)
      memory[3] = 32'b00000010000000001000000000100100; //        and    $s0, $s0, $zero (s0 = 0)
      //memory[4] = 32'b00000000000000000000000000000000; // nop for testing, after testing, we need to stall the sub instruction
     // memory[4] = 32'b00000010001100001000000000100010; //        sub    $s0, $s1, $s0 (s0 = 1)
      memory[4] = 32'b00100000000100000000000000000001; //      addi $s0, $zero, 1 (s0 = 1)
      memory[5] = 32'b00000010000000001000000000100111; //        nor    $s0, $s0, $zero (s0 = -2)
	  memory[6] = 32'b00000010000000001000000000100111;  //		nor	$s0, $s0, $zero (s0 = 1)
	  memory[7] = 32'b00000000000000001000000000100101; //		or	$s0, $zero, $zero (s0 = 0)
	  memory[8] = 32'b00000010001000001000000000100101; //		or	$s0, $s1, $zero (s0 = 1)
	  memory[9] = 32'b00000000000100001000000010000000; //		sll	$s0, $s0, 2 (s0 = 4)
	  memory[10] = 32'b00000010001100001000000000000100; //		sllv	$s0, $s0, $s1 (s0 = 8)*/
		/*Lab 15-17 test case
		memory[0] = 32'b00110100000001000000000000000000;
        memory[1] = 32'b00000000000000000000000000000000;
        memory[2] = 32'b00000000000000000000000000000000;
        memory[3] = 32'b00000000000000000000000000000000;
        memory[4] = 32'b00000000000000000000000000000000;
        memory[5] = 32'b00000000000000000000000000000000;
        memory[6] = 32'b00001000000000000000000000011000;
        memory[7] = 32'b00000000000000000000000000000000;
        memory[8] = 32'b00000000000000000000000000000000;
        memory[9] = 32'b00000000000000000000000000000000;
        memory[10] = 32'b00000000000000000000000000000000;
        memory[11] = 32'b00000000000000000000000000000000;
        memory[12] = 32'b00100000000001000000000000001010;
        memory[13] = 32'b00000000000000000000000000000000;
        memory[14] = 32'b00000000000000000000000000000000;
        memory[15] = 32'b00000000000000000000000000000000;
        memory[16] = 32'b00000000000000000000000000000000;
        memory[17] = 32'b00000000000000000000000000000000;
        memory[18] = 32'b00100000000001000000000000001010;
        memory[19] = 32'b00000000000000000000000000000000;
        memory[20] = 32'b00000000000000000000000000000000;
        memory[21] = 32'b00000000000000000000000000000000;
        memory[22] = 32'b00000000000000000000000000000000;
        memory[23] = 32'b00000000000000000000000000000000;
        memory[24] = 32'b10001100100100000000000000000100;
        memory[25] = 32'b00000000000000000000000000000000;
        memory[26] = 32'b00000000000000000000000000000000;
        memory[27] = 32'b00000000000000000000000000000000;
        memory[28] = 32'b00000000000000000000000000000000;
        memory[29] = 32'b00000000000000000000000000000000;
        memory[30] = 32'b10001100100100000000000000001000;
        memory[31] = 32'b00000000000000000000000000000000;
        memory[32] = 32'b00000000000000000000000000000000;
        memory[33] = 32'b00000000000000000000000000000000;
        memory[34] = 32'b00000000000000000000000000000000;
        memory[35] = 32'b00000000000000000000000000000000;
        memory[36] = 32'b10101100100100000000000000000000;
        memory[37] = 32'b00000000000000000000000000000000;
        memory[38] = 32'b00000000000000000000000000000000;
        memory[39] = 32'b00000000000000000000000000000000;
        memory[40] = 32'b00000000000000000000000000000000;
        memory[41] = 32'b00000000000000000000000000000000;
        memory[42] = 32'b10101100100100000000000000001100;
        memory[43] = 32'b00000000000000000000000000000000;
        memory[44] = 32'b00000000000000000000000000000000;
        memory[45] = 32'b00000000000000000000000000000000;
        memory[46] = 32'b00000000000000000000000000000000;
        memory[47] = 32'b00000000000000000000000000000000;
        memory[48] = 32'b10001100100100010000000000000000;
        memory[49] = 32'b00000000000000000000000000000000;
        memory[50] = 32'b00000000000000000000000000000000;
        memory[51] = 32'b00000000000000000000000000000000;
        memory[52] = 32'b00000000000000000000000000000000;
        memory[53] = 32'b00000000000000000000000000000000;
        memory[54] = 32'b10001100100100100000000000001100;
        memory[55] = 32'b00000000000000000000000000000000;
        memory[56] = 32'b00000000000000000000000000000000;
        memory[57] = 32'b00000000000000000000000000000000;
        memory[58] = 32'b00000000000000000000000000000000;
        memory[59] = 32'b00000000000000000000000000000000;
        memory[60] = 32'b00010010000000000000000000010111;
        memory[61] = 32'b00000000000000000000000000000000;
        memory[62] = 32'b00000000000000000000000000000000;
        memory[63] = 32'b00000000000000000000000000000000;
        memory[64] = 32'b00000000000000000000000000000000;
        memory[65] = 32'b00000000000000000000000000000000;
        memory[66] = 32'b00000010000000001000100000100000;
        memory[67] = 32'b00000000000000000000000000000000;
        memory[68] = 32'b00000000000000000000000000000000;
        memory[69] = 32'b00000000000000000000000000000000;
        memory[70] = 32'b00000000000000000000000000000000;
        memory[71] = 32'b00000000000000000000000000000000;
        memory[72] = 32'b00010010000100010000000000001011;
        memory[73] = 32'b00000000000000000000000000000000;
        memory[74] = 32'b00000000000000000000000000000000;
        memory[75] = 32'b00000000000000000000000000000000;
        memory[76] = 32'b00000000000000000000000000000000;
        memory[77] = 32'b00000000000000000000000000000000;
        memory[78] = 32'b00001000000000000000000101000000;
        memory[79] = 32'b00000000000000000000000000000000;
        memory[80] = 32'b00000000000000000000000000000000;
        memory[81] = 32'b00000000000000000000000000000000;
        memory[82] = 32'b00000000000000000000000000000000;
        memory[83] = 32'b00000000000000000000000000000000;
        memory[84] = 32'b00100000000100001111111111111111;
        memory[85] = 32'b00000000000000000000000000000000;
        memory[86] = 32'b00000000000000000000000000000000;
        memory[87] = 32'b00000000000000000000000000000000;
        memory[88] = 32'b00000000000000000000000000000000;
        memory[89] = 32'b00000000000000000000000000000000;
        memory[90] = 32'b00000110000000011111111110111111;
        memory[91] = 32'b00000000000000000000000000000000;
        memory[92] = 32'b00000000000000000000000000000000;
        memory[93] = 32'b00000000000000000000000000000000;
        memory[94] = 32'b00000000000000000000000000000000;
        memory[95] = 32'b00000000000000000000000000000000;
        memory[96] = 32'b00100010000100000000000000000001;
        memory[97] = 32'b00000000000000000000000000000000;
        memory[98] = 32'b00000000000000000000000000000000;
        memory[99] = 32'b00000000000000000000000000000000;
        memory[100] = 32'b00000000000000000000000000000000;
        memory[101] = 32'b00000000000000000000000000000000;
        memory[102] = 32'b00000110000000010000000000001011;
        memory[103] = 32'b00000000000000000000000000000000;
        memory[104] = 32'b00000000000000000000000000000000;
        memory[105] = 32'b00000000000000000000000000000000;
        memory[106] = 32'b00000000000000000000000000000000;
        memory[107] = 32'b00000000000000000000000000000000;
        memory[108] = 32'b00001000000000000000000101000000;
        memory[109] = 32'b00000000000000000000000000000000;
        memory[110] = 32'b00000000000000000000000000000000;
        memory[111] = 32'b00000000000000000000000000000000;
        memory[112] = 32'b00000000000000000000000000000000;
        memory[113] = 32'b00000000000000000000000000000000;
        memory[114] = 32'b00100000000100001111111111111111;
        memory[115] = 32'b00000000000000000000000000000000;
        memory[116] = 32'b00000000000000000000000000000000;
        memory[117] = 32'b00000000000000000000000000000000;
        memory[118] = 32'b00000000000000000000000000000000;
        memory[119] = 32'b00000000000000000000000000000000;
        memory[120] = 32'b00000000000000000000000000000000;
        memory[121] = 32'b00011110000000000000000000011000;
        memory[122] = 32'b00000000000000000000000000000000;
        memory[123] = 32'b00000000000000000000000000000000;
        memory[124] = 32'b00000000000000000000000000000000;
        memory[125] = 32'b00000000000000000000000000000000;
        memory[126] = 32'b00000000000000000000000000000000;
        memory[127] = 32'b00100000000100000000000000000001;
        memory[128] = 32'b00000000000000000000000000000000;
        memory[129] = 32'b00000000000000000000000000000000;
        memory[130] = 32'b00000000000000000000000000000000;
        memory[131] = 32'b00000000000000000000000000000000;
        memory[132] = 32'b00000000000000000000000000000000;
        memory[133] = 32'b00000000000000000000000000000000;
        memory[134] = 32'b00011110000000000000000000001011;
        memory[135] = 32'b00000000000000000000000000000000;
        memory[136] = 32'b00000000000000000000000000000000;
        memory[137] = 32'b00000000000000000000000000000000;
        memory[138] = 32'b00000000000000000000000000000000;
        memory[139] = 32'b00000000000000000000000000000000;
        memory[140] = 32'b00001000000000000000000101000000;
        memory[141] = 32'b00000000000000000000000000000000;
        memory[142] = 32'b00000000000000000000000000000000;
        memory[143] = 32'b00000000000000000000000000000000;
        memory[144] = 32'b00000000000000000000000000000000;
        memory[145] = 32'b00000000000000000000000000000000;
        memory[146] = 32'b00000110000000000000000000010111;
        memory[147] = 32'b00000000000000000000000000000000;
        memory[148] = 32'b00000000000000000000000000000000;
        memory[149] = 32'b00000000000000000000000000000000;
        memory[150] = 32'b00000000000000000000000000000000;
        memory[151] = 32'b00000000000000000000000000000000;
        memory[152] = 32'b00100000000100001111111111111111;
        memory[153] = 32'b00000000000000000000000000000000;
        memory[154] = 32'b00000000000000000000000000000000;
        memory[155] = 32'b00000000000000000000000000000000;
        memory[156] = 32'b00000000000000000000000000000000;
        memory[157] = 32'b00000000000000000000000000000000;
        memory[158] = 32'b00000110000000000000000000001011;
        memory[159] = 32'b00000000000000000000000000000000;
        memory[160] = 32'b00000000000000000000000000000000;
        memory[161] = 32'b00000000000000000000000000000000;
        memory[162] = 32'b00000000000000000000000000000000;
        memory[163] = 32'b00000000000000000000000000000000;
        memory[164] = 32'b00001000000000000000000101000000;
        memory[165] = 32'b00000000000000000000000000000000;
        memory[166] = 32'b00000000000000000000000000000000;
        memory[167] = 32'b00000000000000000000000000000000;
        memory[168] = 32'b00000000000000000000000000000000;
        memory[169] = 32'b00000000000000000000000000000000;
        memory[170] = 32'b00100000000100011111111111111111;
        memory[171] = 32'b00000000000000000000000000000000;
        memory[172] = 32'b00000000000000000000000000000000;
        memory[173] = 32'b00000000000000000000000000000000;
        memory[174] = 32'b00000000000000000000000000000000;
        memory[175] = 32'b00000000000000000000000000000000;
        memory[176] = 32'b00010110000100010000000000010001;
        memory[177] = 32'b00000000000000000000000000000000;
        memory[178] = 32'b00000000000000000000000000000000;
        memory[179] = 32'b00000000000000000000000000000000;
        memory[180] = 32'b00000000000000000000000000000000;
        memory[181] = 32'b00000000000000000000000000000000;
        memory[182] = 32'b00010110000000000000000000001011;
        memory[183] = 32'b00000000000000000000000000000000;
        memory[184] = 32'b00000000000000000000000000000000;
        memory[185] = 32'b00000000000000000000000000000000;
        memory[186] = 32'b00000000000000000000000000000000;
        memory[187] = 32'b00000000000000000000000000000000;
        memory[188] = 32'b00001000000000000000000101000000;
        memory[189] = 32'b00000000000000000000000000000000;
        memory[190] = 32'b00000000000000000000000000000000;
        memory[191] = 32'b00000000000000000000000000000000;
        memory[192] = 32'b00000000000000000000000000000000;
        memory[193] = 32'b00000000000000000000000000000000;
        memory[194] = 32'b00100000000100000000000010000000;
        memory[195] = 32'b00000000000000000000000000000000;
        memory[196] = 32'b00000000000000000000000000000000;
        memory[197] = 32'b00000000000000000000000000000000;
        memory[198] = 32'b00000000000000000000000000000000;
        memory[199] = 32'b00000000000000000000000000000000;
        memory[200] = 32'b10100000100100000000000000000000;
        memory[201] = 32'b00000000000000000000000000000000;
        memory[202] = 32'b00000000000000000000000000000000;
        memory[203] = 32'b00000000000000000000000000000000;
        memory[204] = 32'b00000000000000000000000000000000;
        memory[205] = 32'b00000000000000000000000000000000;
        memory[206] = 32'b10000000100100000000000000000000;
        memory[207] = 32'b00000000000000000000000000000000;
        memory[208] = 32'b00000000000000000000000000000000;
        memory[209] = 32'b00000000000000000000000000000000;
        memory[210] = 32'b00000000000000000000000000000000;
        memory[211] = 32'b00000000000000000000000000000000;
        memory[212] = 32'b00011010000000000000000000001011;
        memory[213] = 32'b00000000000000000000000000000000;
        memory[214] = 32'b00000000000000000000000000000000;
        memory[215] = 32'b00000000000000000000000000000000;
        memory[216] = 32'b00000000000000000000000000000000;
        memory[217] = 32'b00000000000000000000000000000000;
        memory[218] = 32'b00001000000000000000000101000000;
        memory[219] = 32'b00000000000000000000000000000000;
        memory[220] = 32'b00000000000000000000000000000000;
        memory[221] = 32'b00000000000000000000000000000000;
        memory[222] = 32'b00000000000000000000000000000000;
        memory[223] = 32'b00000000000000000000000000000000;
        memory[224] = 32'b00100000000100001111111111111111;
        memory[225] = 32'b00000000000000000000000000000000;
        memory[226] = 32'b00000000000000000000000000000000;
        memory[227] = 32'b00000000000000000000000000000000;
        memory[228] = 32'b00000000000000000000000000000000;
        memory[229] = 32'b00000000000000000000000000000000;
        memory[230] = 32'b10100100100100000000000000000000;
        memory[231] = 32'b00000000000000000000000000000000;
        memory[232] = 32'b00000000000000000000000000000000;
        memory[233] = 32'b00000000000000000000000000000000;
        memory[234] = 32'b00000000000000000000000000000000;
        memory[235] = 32'b00000000000000000000000000000000;
        memory[236] = 32'b00100000000100000000000000000000;
        memory[237] = 32'b00000000000000000000000000000000;
        memory[238] = 32'b00000000000000000000000000000000;
        memory[239] = 32'b00000000000000000000000000000000;
        memory[240] = 32'b00000000000000000000000000000000;
        memory[241] = 32'b00000000000000000000000000000000;
        memory[242] = 32'b10000100100100000000000000000000;
        memory[243] = 32'b00000000000000000000000000000000;
        memory[244] = 32'b00000000000000000000000000000000;
        memory[245] = 32'b00000000000000000000000000000000;
        memory[246] = 32'b00000000000000000000000000000000;
        memory[247] = 32'b00000000000000000000000000000000;
        memory[248] = 32'b00011010000000000000000000001011;
        memory[249] = 32'b00000000000000000000000000000000;
        memory[250] = 32'b00000000000000000000000000000000;
        memory[251] = 32'b00000000000000000000000000000000;
        memory[252] = 32'b00000000000000000000000000000000;
        memory[253] = 32'b00000000000000000000000000000000;
        memory[254] = 32'b00001000000000000000000101000000;
        memory[255] = 32'b00000000000000000000000000000000;
        memory[256] = 32'b00000000000000000000000000000000;
        memory[257] = 32'b00000000000000000000000000000000;
        memory[258] = 32'b00000000000000000000000000000000;
        memory[259] = 32'b00000000000000000000000000000000;
        memory[260] = 32'b00100000000100001111111111111111;
        memory[261] = 32'b00000000000000000000000000000000;
        memory[262] = 32'b00000000000000000000000000000000;
        memory[263] = 32'b00000000000000000000000000000000;
        memory[264] = 32'b00000000000000000000000000000000;
        memory[265] = 32'b00000000000000000000000000000000;
        memory[266] = 32'b00111100000100000000000000000001;
        memory[267] = 32'b00000000000000000000000000000000;
        memory[268] = 32'b00000000000000000000000000000000;
        memory[269] = 32'b00000000000000000000000000000000;
        memory[270] = 32'b00000000000000000000000000000000;
        memory[271] = 32'b00000000000000000000000000000000;
        memory[272] = 32'b00000110000000010000000000001011;
        memory[273] = 32'b00000000000000000000000000000000;
        memory[274] = 32'b00000000000000000000000000000000;
        memory[275] = 32'b00000000000000000000000000000000;
        memory[276] = 32'b00000000000000000000000000000000;
        memory[277] = 32'b00000000000000000000000000000000;
        memory[278] = 32'b00001000000000000000000101000000;
        memory[279] = 32'b00000000000000000000000000000000;
        memory[280] = 32'b00000000000000000000000000000000;
        memory[281] = 32'b00000000000000000000000000000000;
        memory[282] = 32'b00000000000000000000000000000000;
        memory[283] = 32'b00000000000000000000000000000000;
        memory[284] = 32'b00001000000000000000000100101000;
        memory[285] = 32'b00000000000000000000000000000000;
        memory[286] = 32'b00000000000000000000000000000000;
        memory[287] = 32'b00000000000000000000000000000000;
        memory[288] = 32'b00000000000000000000000000000000;
        memory[289] = 32'b00000000000000000000000000000000;
        memory[290] = 32'b00100010000100001111111111111110;
        memory[291] = 32'b00000000000000000000000000000000;
        memory[292] = 32'b00000000000000000000000000000000;
        memory[293] = 32'b00000000000000000000000000000000;
        memory[294] = 32'b00000000000000000000000000000000;
        memory[295] = 32'b00000000000000000000000000000000;
        memory[296] = 32'b00001100000000000000000100110100;
        memory[297] = 32'b00000000000000000000000000000000;
        memory[298] = 32'b00000000000000000000000000000000;
        memory[299] = 32'b00000000000000000000000000000000;
        memory[300] = 32'b00000000000000000000000000000000;
        memory[301] = 32'b00000000000000000000000000000000;
        memory[302] = 32'b00001000000000000000000000011000;
        memory[303] = 32'b00000000000000000000000000000000;
        memory[304] = 32'b00000000000000000000000000000000;
        memory[305] = 32'b00000000000000000000000000000000;
        memory[306] = 32'b00000000000000000000000000000000;
        memory[307] = 32'b00000000000000000000000000000000;
        memory[308] = 32'b00000011111000000000000000001000;
        memory[309] = 32'b00000000000000000000000000000000;
        memory[310] = 32'b00000000000000000000000000000000;
        memory[311] = 32'b00000000000000000000000000000000;
        memory[312] = 32'b00000000000000000000000000000000;
        memory[313] = 32'b00000000000000000000000000000000;
        memory[314] = 32'b00001000000000000000000101000000;
        memory[315] = 32'b00000000000000000000000000000000;
        memory[316] = 32'b00000000000000000000000000000000;
        memory[317] = 32'b00000000000000000000000000000000;
        memory[318] = 32'b00000000000000000000000000000000;
        memory[319] = 32'b00000000000000000000000000000000;
        memory[320] = 32'b00000000000000000000000000001000;
        memory[321] = 32'b00000000000000000000000000000000;
        memory[322] = 32'b00000000000000000000000000000000;
        memory[323] = 32'b00000000000000000000000000000000;
        memory[324] = 32'b00000000000000000000000000000000;
        memory[325] = 32'b00000000000000000000000000000000;
        memory[326] = 32'b00110100000000100000000000001010;
        memory[327] = 32'b00000000000000000000000000000000;
        memory[328] = 32'b00000000000000000000000000000000;
        memory[329] = 32'b00000000000000000000000000000000;
        memory[330] = 32'b00000000000000000000000000000000;
        memory[331] = 32'b00000000000000000000000000000000;
        memory[332] = 32'b00000000000000000000000000000000;
        memory[333] = 32'b00000000000000000000000000000000;
        memory[334] = 32'b00000000000000000000000000000000;
        memory[335] = 32'b00000000000000000000000000000000;
        memory[336] = 32'b00000000000000000000000000000000;
        memory[337] = 32'b00000000000000000000000000000000;*/

	end
	
	always@(*) begin
	   Instruction <= memory[Address[11:2]];
	end
	
endmodule
